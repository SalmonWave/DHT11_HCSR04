`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: T.Y JANG
// 
// Create Date: 12/11/2024 01:50:25 PM
// Design Name: 
// Module Name: COUNTER FOR CLOCK
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module counter_6000_clock (
    input                       clk,
    input                       i_tick,
    input                       reset,
    output [$clog2(11600) - 1:0] o_bcd
);

////////////////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////  WIRE & REG   ////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////

    reg [$clog2(6_000)-1:0] count, count_next;


////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////  MODULE Logic   ////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////

    always @(posedge clk, posedge reset) begin
        if (reset) begin
            count <= 0;
        end else begin
            count <= count_next;
        end
    end

    always @(*) begin

        count_next = count;


        if (i_tick) begin
            if (count == 6_000) begin
                count_next = 0;
            end else begin
                count_next = count + 1;
            end
        end

    end

    assign o_bcd = count;

endmodule


module tick_10ms_clock (
    input clk,
    input reset,
    output reg tick_100hz
);


////////////////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////  WIRE & REG   ////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////

    reg [$clog2(1_000_000)-1:0] r_counter;  


////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////  MODULE Logic   ////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////


    always @(posedge clk, posedge reset) begin


        if (reset) begin
            r_counter  <= 0;
            tick_100hz <= 0;


        end else begin
            if (r_counter == 1_000_000) begin
                r_counter  <= 0;
                tick_100hz <= 1'b1;
            end else begin
                r_counter  <= r_counter + 1;
                tick_100hz <= 1'b0;
            end
        end
    end

endmodule











module counter_minute_count_clock (
    input clk,
    input i_tick,
    input reset,
    output [$clog2(11600) - 1:0] o_bcd
);

 ////////////////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////  WIRE & REG   ////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////

    reg [$clog2(60)-1:0] count, count_next;
    reg [$clog2(1_000)-1:0] minute_counter, minute_counter_next;


////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////  MODULE Logic   ////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////

    always @(posedge clk, posedge reset) begin
        if (reset) begin
            count <= 0;
            minute_counter <= 0;
        end else begin
            count <= count_next;
            minute_counter <= minute_counter_next;
        end
    end


    always @(*) begin

        count_next = count;
        minute_counter_next = minute_counter;

        if (i_tick) begin
            if (count == 59) begin
                count_next = 0;
                minute_counter_next = minute_counter + 1;
                if(minute_counter == 1_000) begin
                    minute_counter_next = 0;
                end

            end else begin
                count_next = count + 1;
            end
        end
    end
    
    assign o_bcd = minute_counter;

endmodule


module tick_1Hz_clock (
    input clk,
    input reset,
    output reg tick_1hz
);

////////////////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////  WIRE & REG   ////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////

    reg [$clog2(100_000_000)-1:0] r_counter;


////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////  MODULE Logic   ////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////

    always @(posedge clk, posedge reset) begin

        if (reset) begin
            r_counter  <= 0;
            tick_1hz <= 0;


        end else begin
            if (r_counter == 100_000_000) begin
                r_counter  <= 0;
                tick_1hz <= 1'b1;
            end else begin
                r_counter  <= r_counter + 1;
                tick_1hz <= 1'b0;
            end
        end
    end


endmodule
